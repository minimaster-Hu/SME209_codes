`timescale 1ns / 1ps

module mem(
    input clk,
    input [7:0] addr,
    output reg [31:0] data
);

// TODO  
    
endmodule
